module mem
(
    input  logic in, 
    output logic out
);

assign out = in;

logic [31:0] mem [9999:0];

endmodule