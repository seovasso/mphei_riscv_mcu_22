module mpei_rv_top (
);
endmodule 
